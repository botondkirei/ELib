��l i b r a r y   I E E E ;  
 u s e   I E E E . s t d _ l o g i c _ 1 1 6 4 . a l l ;  
  
  
 p a c k a g e   P A E C o r e   i s    
  
 	  
 	 t y p e   A t y p e   i s   p r o t e c t e d  
 	 	 p r o c e d u r e   a d d A r e a ( i n c r e m e n t   :   r e a l   ; c o n s t a n t   D o m a i n   :   i n t e g e r   )   ;  
 	 	 p r o c e d u r e   r e p o r t A r e a ( c o n s t a n t   D o m a i n   :   i n t e g e r ) ;  
 	 e n d   p r o t e c t e d   A t y p e ;  
 	  
 	 s h a r e d   v a r i a b l e   A M   :   A t y p e ;    
  
 	 t y p e   P t y p e   i s   p r o t e c t e d  
 	 	 p r o c e d u r e   a d d L e a c k a g e ( c o n s t a n t   p l e a c k :   r e a l   ;   c o n s t a n t   D o m a i n   :   i n t e g e r ) ;  
 	 	 p r o c e d u r e   i n c ( v a r i a b l e   i n c r e m e n t   :   r e a l ;   c o n s t a n t   D o m a i n   :   i n t e g e r ) ;  
 	 	 p r o c e d u r e   r e p o r t P o w e r ( c o n s t a n t   D o m a i n :   i n t e g e r ) ;  
 	 	 p r o c e d u r e   r e s e t P o w e r ( c o n s t a n t   D o m a i n :   i n t e g e r ) ;  
 	 	 i m p u r e   f u n c t i o n   g e t P o w e r ( c o n s t a n t   D o m a i n   :   i n t e g e r )   r e t u r n   r e a l ;  
 	 	 p r o c e d u r e   m o n i t o r I n p u t ( s i g n a l   i n p u t :   s t d _ l o g i c ;   c o n s t a n t   C   :   r e a l   ;   s i g n a l   s u p p l y   :   r e a l ;   c o n s t a n t   D o m a i n   :   i n t e g e r )   ; 	  
 	 	 p r o c e d u r e   m o n i t o r I n p u t ( s i g n a l   i n p u t :   s t d _ l o g i c _ v e c t o r ;   c o n s t a n t   C   :   r e a l   ;   s i g n a l   s u p p l y   :   r e a l ;   c o n s t a n t   D o m a i n   :   i n t e g e r )   ; 	  
 	 e n d   p r o t e c t e d   P t y p e ;  
 	  
 	 s h a r e d   v a r i a b l e   P M :   P t y p e ;  
 	  
 	 t y p e   r e a l _ a r r a y   i s   a r r a y   ( 1   t o   1 6 )   o f   r e a l ;  
 	  
 e n d   P A E C o r e ;  
  
 p a c k a g e   b o d y     P A E C o r e   i s  
  
 	 t y p e   P t y p e   i s   p r o t e c t e d   b o d y  
 	  
 	 	 v a r i a b l e   s o c k e t   :   r e a l _ a r r a y   : =   ( o t h e r s   = >   0 . 0 ) ;  
 	 	 v a r i a b l e   l e a c k   :   r e a l _ a r r a y   : =   ( o t h e r s   = >   0 . 0 ) ;  
 	 	  
 	 	 p r o c e d u r e   a d d L e a c k a g e ( c o n s t a n t   p l e a c k :   r e a l   ;   c o n s t a n t   D o m a i n   :   i n t e g e r )   i s  
 	 	 b e g i n  
 	 	 	 l e a c k ( D o m a i n )   : =   l e a c k ( D o m a i n )   +   p l e a c k ;  
 	 	 e n d   p r o c e d u r e ;  
  
 	 	 p r o c e d u r e   i n c   ( v a r i a b l e   i n c r e m e n t   :   r e a l ;   c o n s t a n t   D o m a i n   :   i n t e g e r )   i s  
 	 	 b e g i n  
 	 	 	 s o c k e t ( D o m a i n )   : =   s o c k e t ( D o m a i n )   +   i n c r e m e n t ;  
 	 	 e n d   p r o c e d u r e ;  
 	 	  
 	 	 p r o c e d u r e   r e p o r t P o w e r ( c o n s t a n t   D o m a i n :   i n t e g e r )   i s  
 	 	 b e g i n  
 	 	 	 r e p o r t   " D o m a i n   "   &   i n t e g e r ' i m a g e   ( D o m a i n )   &   "   d y n a m i c   p o w e r   ( J o u l e ) :   "   &   r e a l ' i m a g e ( s o c k e t ( D o m a i n ) ) ;  
 	 	 	 r e p o r t   " D o m a i n   "   &   i n t e g e r ' i m a g e   ( D o m a i n )   &   "   l e a c k a g e   p o w e r   ( n W ) :   "   &   r e a l ' i m a g e ( l e a c k ( D o m a i n ) ) ;  
 	 	 e n d   p r o c e d u r e ;  
 	 	  
 	 	 p r o c e d u r e   r e s e t P o w e r ( c o n s t a n t   D o m a i n :   i n t e g e r )   i s  
 	 	 b e g i n  
 	 	 	 s o c k e t ( D o m a i n )   : =   0 . 0 ;  
 	 	 e n d   p r o c e d u r e ;  
 	 	  
 	 	 i m p u r e   f u n c t i o n   g e t P o w e r ( c o n s t a n t   D o m a i n   :   i n t e g e r )   r e t u r n   r e a l   i s  
 	 	 b e g i n  
 	 	 	 r e t u r n   s o c k e t ( D o m a i n ) ;  
 	 	 e n d   f u n c t i o n ;  
 	 	  
 	 	 p r o c e d u r e   m o n i t o r I n p u t ( s i g n a l   i n p u t :   s t d _ l o g i c ;   c o n s t a n t   C   :   r e a l   ;   s i g n a l   s u p p l y   :   r e a l ;   c o n s t a n t   D o m a i n   :   i n t e g e r )   i s  
 	 	 	 v a r i a b l e   i n c r e m e n t   :   r e a l   : =   1 . 0 ;  
 	 	 b e g i n  
 	 	 	 i n c r e m e n t   : =   s u p p l y * s u p p l y * C   /   2 . 0 ;  
 	 	 	 i f   i n p u t ' e v e n t   t h e n  
 	 	 	 	 i n c ( i n c r e m e n t , D o m a i n ) ;  
 	 	 	 e n d   i f ;  
 	 	 e n d   p r o c e d u r e ;  
  
 	 	 p r o c e d u r e   m o n i t o r I n p u t ( s i g n a l   i n p u t :   s t d _ l o g i c _ v e c t o r ;   c o n s t a n t   C   :   r e a l   ;   s i g n a l   s u p p l y   :   r e a l ;   c o n s t a n t   D o m a i n   :   i n t e g e r )   i s  
 	 	 	 v a r i a b l e   i n c r e m e n t   :   r e a l   : =   1 . 0 ;  
 	 	 b e g i n  
 	 	 	 i n c r e m e n t   : =   s u p p l y * s u p p l y * C   /   2 . 0 ;  
 	 	 	 f o r   i   i n   0   t o   i n p u t ' l e n g t h   -   1   l o o p  
 	 	 	 	 i f   i n p u t ( i ) ' e v e n t   t h e n  
 	 	 	 	 	 i n c ( i n c r e m e n t , D o m a i n ) ;  
 	 	 	 	 e n d   i f ;  
 	 	 	 e n d   l o o p ;  
 	 	 e n d   p r o c e d u r e ;  
 	 	 	 	  
 	 e n d   p r o t e c t e d   b o d y   P t y p e ;  
 	  
 	 t y p e   A t y p e   i s   p r o t e c t e d   b o d y  
 	  
 	 	 v a r i a b l e   t o t a l A r e a   :   r e a l _ a r r a y   : =   ( o t h e r s   = >   0 . 0 ) ;  
 	  
 	 	 p r o c e d u r e   a d d A r e a ( i n c r e m e n t   :   r e a l   ;   c o n s t a n t   D o m a i n   :   i n t e g e r )   i s  
 	 	 b e g i n  
 	 	 	 t o t a l A r e a ( D o m a i n )   : =   t o t a l A r e a ( D o m a i n )   +   i n c r e m e n t ;  
 	 	 e n d   p r o c e d u r e ;  
 	 	  
 	 	 p r o c e d u r e   r e p o r t A r e a ( c o n s t a n t   D o m a i n   :   i n t e g e r )   i s  
 	 	 b e g i n  
 	 	 	 r e p o r t   " D o m a i n   "   &   i n t e g e r ' i m a g e   ( D o m a i n )   &   "   a r e a :   "   &   r e a l ' i m a g e ( t o t a l A r e a ( D o m a i n ) ) ;  
 	 	 e n d   p r o c e d u r e ;  
 	 	  
 	 e n d   p r o t e c t e d   b o d y   A t y p e ;  
 	  
  
 	  
 e n d   p a c k a g e   b o d y ;  
 