library ieee;
use ieee.std_logic_vector.all;

package sxlib is

  component 
  end compnent
  
end package;

package body sxlib is

end package body;
